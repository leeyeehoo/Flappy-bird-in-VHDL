LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY BIRD IS
	PORT(
		 CLK_OUT:OUT STD_LOGIC;
		 CLK_IN:IN STD_LOGIC;		 
		 CONTROL_BTN:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 CONTROL_BTN2:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 RESET_BTN:IN STD_LOGIC;
	     R_COL:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 ROW:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 G_COL:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 NUM:OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
		 CAT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		 SPEED_BTN:IN STD_LOGIC;
		 MODE_BTN:IN STD_LOGIC;
		 MODE_LIGHT:OUT STD_LOGIC;
		 BEEP:OUT STD_LOGIC;
		 RW,EN,RS:OUT STD_LOGIC;
         QDATA:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
		 );
END BIRD;
ARCHITECTURE IGNIGHT OF BIRD IS
	SIGNAL CLK:STD_LOGIC;
	SIGNAL TMP_MAIN:INTEGER RANGE 0 TO 24999;
	SIGNAL TMP:INTEGER RANGE 0 TO 7;
	SIGNAL TMP_DOUBLE:INTEGER RANGE 0 TO 15;
	SIGNAL COUNT:INTEGER RANGE 0 TO 1;
	SIGNAL DTMP:INTEGER RANGE 0 TO 499;
	SIGNAL TMP_SOUND:INTEGER RANGE 0 TO 6249999;
	SIGNAL CLKTMP:STD_LOGIC;
	SIGNAL CLK_SOUND:STD_LOGIC;
	SIGNAL STMP:INTEGER RANGE 0 TO 49;
	SIGNAL CLK_ANTISHAKE:STD_LOGIC;
	SIGNAL CLK_BEEP:STD_LOGIC;
	SIGNAL MOVE:INTEGER RANGE 0 TO 33;
	SIGNAL MOVE_FLAG:INTEGER RANGE 0 TO 11;
	SIGNAL POSITION:INTEGER RANGE 0 TO 7;
	SIGNAL POSITION2:INTEGER RANGE 0 TO 7;
	SIGNAL FAIL_FLAG:INTEGER RANGE 0 TO 1;
	SIGNAL FAIL_FLAG2:INTEGER RANGE 0 TO 1;
	SIGNAL RESET:INTEGER RANGE 0 TO 1;
	SIGNAL CAT_TMP:INTEGER RANGE 0 TO 1;
	SIGNAL RAM:STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL FEEDBACK:STD_LOGIC;
	SIGNAL TUBE1:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TUBE2:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TUBE3:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TUBE4:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TUBE5:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TUBE6:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TUBE0:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP1:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP2:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP3:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP4:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP5:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP6:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP7:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL G_COL_TMP8:STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL LINE1:INTEGER RANGE 0 TO 6;
	SIGNAL LINE2:INTEGER RANGE 0 TO 6;
	SIGNAL LINE3:INTEGER RANGE 0 TO 6;
	SIGNAL NUM_TMP1:STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL NUM_TMP2:STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL MODE:INTEGER RANGE 0 TO 1;
	SIGNAL MODE_TMP:INTEGER RANGE 0 TO 1;
	SIGNAL WIN:INTEGER RANGE 0 TO 2;
	SIGNAL SELECTION:INTEGER RANGE 0 TO 127;
	SIGNAL TUNE:INTEGER RANGE 0 TO 75758;
	SIGNAL CNT:INTEGER RANGE 0 TO 75758;
	CONSTANT MI:INTEGER:= 75758;------330 75758
	CONSTANT FA:INTEGER:= 67568;------370 67568
	CONSTANT SO:INTEGER:= 63776;------392 63776
	CONSTANT LA:INTEGER:= 56818;------440 56818
	CONSTANT XI:INTEGER:= 50607;------494 50607
	CONSTANT DO_HIGH:INTEGER:= 47801;------523 47801
	CONSTANT DO_HIGH2:INTEGER:= 45126;------554 45126
	CONSTANT RE_HIGH:INTEGER:= 42589;------587 42589
	CONSTANT MI_HIGH:INTEGER:=37936;------659 37936
	BEGIN
	RW<='0';
    EN<=CLK;
    P0:PROCESS(CLK_IN)
		BEGIN
		IF CLK_IN'EVENT AND CLK_IN='1' THEN
			IF TMP_MAIN=24999 THEN
				TMP_MAIN<=0;
				CLK<=NOT CLK;
			ELSE
				TMP_MAIN<=TMP_MAIN+1;
			END IF;
		END IF;
		END PROCESS;		
-------------------------------------------------FENPIN1
	P1:PROCESS(CLK,SPEED_BTN)
	BEGIN
		IF CLK'EVENT AND CLK='1' THEN
		IF SPEED_BTN='1' THEN
			IF DTMP=499 THEN
				DTMP<=0;
				CLKTMP<=NOT CLKTMP;
			ELSE
				DTMP<=DTMP+1;
			END IF;
		ELSIF SPEED_BTN='0' THEN
			IF DTMP=249 THEN
				DTMP<=0;
				CLKTMP<=NOT CLKTMP;
			ELSIF DTMP=499 THEN
				DTMP<=250;
				CLKTMP<=NOT CLKTMP;
			ELSE
				DTMP<=DTMP+1;
			END IF;
		END IF;
		END IF;		
	CLK_OUT<=CLKTMP;
	END PROCESS;
-------------------------------------------------SAOMIAO
	P2:PROCESS(DTMP)
	BEGIN
		TMP<=DTMP MOD 8;
	END PROCESS;
	P3:PROCESS(TMP)
	BEGIN 
		CASE TMP IS
			WHEN 0=>ROW<="11111110";
			WHEN 1=>ROW<="11111101";
			WHEN 2=>ROW<="11111011";
			WHEN 3=>ROW<="11110111";
			WHEN 4=>ROW<="11101111";
			WHEN 5=>ROW<="11011111";
			WHEN 6=>ROW<="10111111";
			WHEN 7=>ROW<="01111111";
		END CASE;
	END PROCESS;
-------------------------------------------------MOVE
	P4:PROCESS(CLKTMP,FAIL_FLAG,FAIL_FLAG2,RESET)
	BEGIN
		IF CLKTMP'EVENT AND CLKTMP='1' THEN
			IF MOVE=32 OR MOVE=33 THEN
				MOVE<=MOVE;			
			ELSE 
				IF FAIL_FLAG=0 AND FAIL_FLAG2=0 THEN
				MOVE<=MOVE+1;
				ELSIF FAIL_FLAG=1 OR FAIL_FLAG2=1 THEN
					IF FAIL_FLAG=1 AND FAIL_FLAG2=1 THEN
						WIN<=0;
					ELSIF FAIL_FLAG=1 AND FAIL_FLAG2=0 THEN
						WIN<=1;
					ELSE
						WIN<=2;
					END IF;
				MOVE<=33;
				END IF;
			END IF;					
		END IF;
		
		IF RESET=1 THEN
		MOVE<=0;
		END IF;
		IF MODE_TMP=1 THEN
			MOVE<=0;
		END IF;
	END PROCESS;
	P5:PROCESS(CLKTMP,MOVE)
	BEGIN
		IF CLKTMP'EVENT AND CLKTMP='1' THEN
			IF MOVE=0 OR MOVE =1  THEN
				COUNT<=0;
			ELSE
				IF COUNT=0 THEN
					COUNT<=COUNT+1;
				ELSE COUNT<=0;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	P6:PROCESS(CLKTMP,RAM,COUNT)
	BEGIN
		IF CLKTMP'EVENT AND CLKTMP='1' THEN			
			TUBE1<="00011111";
			TUBE2<="10001111";
			TUBE3<="11000111";
			TUBE4<="11100011";
			TUBE5<="11110001";
			TUBE6<="11111000";
			TUBE0<="00000000";
			IF MOVE=0 OR MOVE=1 OR MOVE=32 OR MOVE=33 THEN
					G_COL_TMP1<="00000000";
					G_COL_TMP2<="00000000";
					G_COL_TMP3<="00000000";
					G_COL_TMP4<="00000000";
					G_COL_TMP5<="00000000";
					G_COL_TMP6<="00000000";
					G_COL_TMP7<="00000000";
					G_COL_TMP8<="00000000";
					LINE1<=0;
					LINE2<=0;
					LINE3<=0;
			ELSE
			IF COUNT=1 THEN
				IF RAM="0000" OR RAM="0001" OR RAM="0010" THEN
					G_COL_TMP1<=TUBE1(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE1(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE1(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE1(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE1(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE1(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE1(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE1(0)&G_COL_TMP8(7 DOWNTO 1);
					LINE3<=LINE2;
					LINE2<=LINE1;
					LINE1<=1;
				ELSIF RAM="0011" OR RAM="0100" OR RAM="0101" THEN
					G_COL_TMP1<=TUBE2(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE2(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE2(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE2(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE2(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE2(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE2(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE2(0)&G_COL_TMP8(7 DOWNTO 1);
					LINE3<=LINE2;
					LINE2<=LINE1;
					LINE1<=2;
				ELSIF RAM="0110" OR RAM="0111" OR RAM="1000" THEN
					G_COL_TMP1<=TUBE3(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE3(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE3(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE3(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE3(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE3(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE3(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE3(0)&G_COL_TMP8(7 DOWNTO 1);
					LINE3<=LINE2;
					LINE2<=LINE1;
					LINE1<=3;
				ELSIF RAM="1001" OR RAM="1010"  THEN
					G_COL_TMP1<=TUBE4(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE4(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE4(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE4(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE4(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE4(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE4(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE4(0)&G_COL_TMP8(7 DOWNTO 1);
					LINE3<=LINE2;
					LINE2<=LINE1;
					LINE1<=4;
				ELSIF RAM="1011" OR RAM="1100"  THEN
					G_COL_TMP1<=TUBE5(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE5(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE5(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE5(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE5(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE5(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE5(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE5(0)&G_COL_TMP8(7 DOWNTO 1);
					LINE3<=LINE2;
					LINE2<=LINE1;
					LINE1<=5;
				ELSIF RAM="1101" OR RAM="1110" OR RAM="1111" THEN
					G_COL_TMP1<=TUBE6(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE6(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE6(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE6(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE6(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE6(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE6(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE6(0)&G_COL_TMP8(7 DOWNTO 1);
					LINE3<=LINE2;
					LINE2<=LINE1;
					LINE1<=6;
				
				END IF;
			ELSE
					G_COL_TMP1<=TUBE0(7)&G_COL_TMP1(7 DOWNTO 1);
					G_COL_TMP2<=TUBE0(6)&G_COL_TMP2(7 DOWNTO 1);
					G_COL_TMP3<=TUBE0(5)&G_COL_TMP3(7 DOWNTO 1);
					G_COL_TMP4<=TUBE0(4)&G_COL_TMP4(7 DOWNTO 1);
					G_COL_TMP5<=TUBE0(3)&G_COL_TMP5(7 DOWNTO 1);
					G_COL_TMP6<=TUBE0(2)&G_COL_TMP6(7 DOWNTO 1);
					G_COL_TMP7<=TUBE0(1)&G_COL_TMP7(7 DOWNTO 1);
					G_COL_TMP8<=TUBE0(0)&G_COL_TMP8(7 DOWNTO 1);
			END IF;
		END IF;
		END IF;
	END PROCESS;
	P7:PROCESS(LINE3,COUNT,MODE,POSITION,POSITION2)
	BEGIN
	IF MODE=0 THEN
		IF COUNT=1 THEN
			CASE LINE3 IS
				WHEN 0=>
					FAIL_FLAG<=0;
				WHEN 6=>
					IF POSITION=0 OR POSITION=1 OR POSITION=2 OR  POSITION=3 OR POSITION=4 THEN 
					FAIL_FLAG<=1;					
					ELSE 
					FAIL_FLAG<=0;	
					END IF;								
				WHEN 5=>
					IF POSITION=0 OR POSITION=1 OR POSITION=2 OR  POSITION=3 OR POSITION=7 THEN 
					FAIL_FLAG<=1;					
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
				WHEN 4=>
					IF POSITION=0 OR POSITION=1 OR POSITION=2 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;					
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
				WHEN 3=>
					IF POSITION=0 OR POSITION=1 OR POSITION=5 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;					
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
				WHEN 2=>
					IF POSITION=0 OR POSITION=4 OR POSITION=5 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;					
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
				WHEN 1=>
					IF POSITION=3 OR POSITION=4 OR POSITION=5 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;					
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
			END CASE;
		ELSE
			FAIL_FLAG<=0;
		END IF;
	ELSE
		IF COUNT=1 THEN
			CASE LINE3 IS
				WHEN 0=>
					FAIL_FLAG<=0;
					FAIL_FLAG2<=0;
				WHEN 6=>
					IF POSITION=0 OR POSITION=1 OR POSITION=2 OR  POSITION=3 OR POSITION=4 THEN 
					FAIL_FLAG<=1;
					ELSE 
					FAIL_FLAG<=0;	
					END IF;				
					IF POSITION2=0 OR POSITION2=1 OR POSITION2=2 OR  POSITION2=3 OR POSITION2=4 THEN 
					FAIL_FLAG2<=1;
					ELSE 
					FAIL_FLAG2<=0;	
					END IF;				
				WHEN 5=>
					IF POSITION=0 OR POSITION=1 OR POSITION=2 OR  POSITION=3 OR POSITION=7 THEN 
					FAIL_FLAG<=1;
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
					IF POSITION2=0 OR POSITION2=1 OR POSITION2=2 OR  POSITION2=3 OR POSITION2=7 THEN 
					FAIL_FLAG2<=1;
					ELSE 
					FAIL_FLAG2<=0;
					END IF;						
				WHEN 4=>
					IF POSITION=0 OR POSITION=1 OR POSITION=2 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
					IF POSITION2=0 OR POSITION2=1 OR POSITION2=2 OR  POSITION2=6 OR POSITION2=7 THEN 
					FAIL_FLAG2<=1;
					ELSE 
					FAIL_FLAG2<=0;
					END IF;						
				WHEN 3=>
					IF POSITION=0 OR POSITION=1 OR POSITION=5 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;	
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
					IF POSITION2=0 OR POSITION2=1 OR POSITION2=5 OR  POSITION2=6 OR POSITION2=7 THEN 
					FAIL_FLAG2<=1;	
					ELSE 
					FAIL_FLAG2<=0;
					END IF;						
				WHEN 2=>
					IF POSITION=0 OR POSITION=4 OR POSITION=5 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;	
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
					IF POSITION2=0 OR POSITION2=4 OR POSITION2=5 OR  POSITION2=6 OR POSITION2=7 THEN 
					FAIL_FLAG2<=1;	
					ELSE 
					FAIL_FLAG2<=0;
					END IF;						
				WHEN 1=>
					IF POSITION=3 OR POSITION=4 OR POSITION=5 OR  POSITION=6 OR POSITION=7 THEN 
					FAIL_FLAG<=1;	
					ELSE 
					FAIL_FLAG<=0;
					END IF;	
					IF POSITION2=3 OR POSITION2=4 OR POSITION2=5 OR  POSITION2=6 OR POSITION2=7 THEN 
					FAIL_FLAG2<=1;			
					ELSE 
					FAIL_FLAG2<=0;
					END IF;						
			END CASE;
		ELSE
			FAIL_FLAG<=0;
			FAIL_FLAG2<=0;
		END IF;
	END IF;
	END PROCESS;
	P8:PROCESS(TMP, MOVE, G_COL_TMP1, G_COL_TMP2, G_COL_TMP3, G_COL_TMP4, G_COL_TMP5, G_COL_TMP6, G_COL_TMP7, G_COL_TMP8)
	BEGIN		
		IF MOVE=0 OR MOVE=1 OR MOVE=2 OR MOVE=32 OR MOVE=33 THEN
				CASE TMP IS
					WHEN 0=>G_COL<="00000000";
					WHEN 1=>G_COL<="00000000";
					WHEN 2=>G_COL<="00000000";
					WHEN 3=>G_COL<="00000000";
					WHEN 4=>G_COL<="00000000";
					WHEN 5=>G_COL<="00000000";
					WHEN 6=>G_COL<="00000000";
					WHEN 7=>G_COL<="00000000";
				END CASE;
		ELSE
				CASE TMP IS
					WHEN 0=>G_COL<=G_COL_TMP1;
					WHEN 1=>G_COL<=G_COL_TMP2;
					WHEN 2=>G_COL<=G_COL_TMP3;
					WHEN 3=>G_COL<=G_COL_TMP4;
					WHEN 4=>G_COL<=G_COL_TMP5;
					WHEN 5=>G_COL<=G_COL_TMP6;
					WHEN 6=>G_COL<=G_COL_TMP7;
					WHEN 7=>G_COL<=G_COL_TMP8;
				END CASE;
		END IF;
	END PROCESS;
-------------------------------------------------XIAONIAO
	P9:PROCESS(CLK)
	BEGIN
	IF CLK'EVENT AND CLK='1' THEN
			IF STMP=49 THEN
				STMP<=0;
				CLK_ANTISHAKE<=NOT CLK_ANTISHAKE;
			ELSE
			STMP<=STMP+1;
			END IF;
			END IF;
	END PROCESS;
	P10:PROCESS(CONTROL_BTN,CLK_ANTISHAKE)
	BEGIN
	IF CLK_ANTISHAKE'EVENT AND CLK_ANTISHAKE='1' AND FAIL_FLAG=0 THEN
		CASE CONTROL_BTN IS
					WHEN "00"=>POSITION<=POSITION;
					WHEN "01"=>
						IF POSITION<7 THEN
							POSITION<=POSITION+1;
						END IF;
						
					WHEN "10"=>
						IF POSITION>0 THEN
							POSITION<=POSITION-1;
						END IF;
					WHEN "11"=>POSITION<=POSITION;
		END CASE;
	END IF;
	END PROCESS;
	P11:PROCESS(POSITION,MOVE,TMP,TMP_DOUBLE,WIN,POSITION2)
	BEGIN
	IF MODE=0 THEN
		IF MOVE/=32 AND MOVE/=33 AND MOVE/=0 AND MOVE/=1 AND MOVE/=2 THEN 
			CASE POSITION IS
			WHEN 0=>CASE TMP IS
					WHEN 0=>R_COL<="00000100";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000000";
				END CASE;
			WHEN 1=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000100";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000000";
				END CASE;
			WHEN 2=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000100";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000000";	
				END CASE;
			WHEN 3=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000100";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000000";	
				END CASE;
			WHEN 4=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000100";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000000";	
				END CASE;
			WHEN 5=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000100";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000000";	
				END CASE;
			WHEN 6=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000100";
					WHEN 7=>R_COL<="00000000";
				END CASE;	
			WHEN 7=>CASE TMP IS
					WHEN 0=>R_COL<="00000000";
					WHEN 1=>R_COL<="00000000";
					WHEN 2=>R_COL<="00000000";
					WHEN 3=>R_COL<="00000000";
					WHEN 4=>R_COL<="00000000";
					WHEN 5=>R_COL<="00000000";
					WHEN 6=>R_COL<="00000000";
					WHEN 7=>R_COL<="00000100";
				END CASE;		
			END CASE;
		ELSIF MOVE=32 THEN
			CASE TMP IS
					WHEN 0=>R_COL<="00011000";
					WHEN 1=>R_COL<="00011000";
					WHEN 2=>R_COL<="00100100";
					WHEN 3=>R_COL<="00100100";
					WHEN 4=>R_COL<="01000010";
					WHEN 5=>R_COL<="01000010";
					WHEN 6=>R_COL<="10000001";
					WHEN 7=>R_COL<="10000001";
				END CASE;
		ELSIF MOVE=33 THEN
			CASE TMP IS
					WHEN 0=>R_COL<="10000001";
					WHEN 1=>R_COL<="01000010";
					WHEN 2=>R_COL<="00100100";
					WHEN 3=>R_COL<="00011000";
					WHEN 4=>R_COL<="00011000";
					WHEN 5=>R_COL<="00100100";
					WHEN 6=>R_COL<="01000010";
					WHEN 7=>R_COL<="10000001";
				END CASE;
		ELSIF MOVE=0 THEN
			CASE TMP IS
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="00011000";
					WHEN 2=>R_COL<="00011000";
					WHEN 3=>R_COL<="00011000";
					WHEN 4=>R_COL<="00011000";
					WHEN 5=>R_COL<="00011000";
					WHEN 6=>R_COL<="00011110";
					WHEN 7=>R_COL<="00011000";
				END CASE;
		ELSIF MOVE=1 THEN
			CASE TMP IS
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="00000011";
					WHEN 2=>R_COL<="00000011";
					WHEN 3=>R_COL<="00000011";
					WHEN 4=>R_COL<="11111111";
					WHEN 5=>R_COL<="11000000";
					WHEN 6=>R_COL<="11000000";
					WHEN 7=>R_COL<="11111111";
				END CASE;
		ELSIF MOVE=2 THEN
			CASE TMP IS
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="10000000";
					WHEN 2=>R_COL<="10000000";
					WHEN 3=>R_COL<="10000000";
					WHEN 4=>R_COL<="11111100";
					WHEN 5=>R_COL<="10000000";
					WHEN 6=>R_COL<="10000000";
					WHEN 7=>R_COL<="11111111";
				END CASE;	
		END IF;
	ELSE
		IF MOVE/=32 AND MOVE/=33 AND MOVE/=0 AND MOVE/=1 AND MOVE/=2 THEN 
			CASE POSITION IS
			WHEN 0=>IF TMP_DOUBLE=0 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;
			WHEN 1=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;
			WHEN 2=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;
			WHEN 3=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;
			WHEN 4=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;
			WHEN 5=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;
			WHEN 6=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000000";
					END IF;	
			WHEN 7=>IF TMP_DOUBLE=0 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=1 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=2 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=3 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=4 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=5 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=6 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=7 THEN R_COL<="00000100";
					END IF;		
			END CASE;
			CASE POSITION2 IS
			WHEN 0=>IF TMP_DOUBLE=8 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;
			WHEN 1=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;
			WHEN 2=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;
			WHEN 3=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;
			WHEN 4=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;
			WHEN 5=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;
			WHEN 6=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000100";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000000";
					END IF;	
			WHEN 7=>IF TMP_DOUBLE=8 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=9 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=10 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=11 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=12 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=13 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=14 THEN R_COL<="00000000";
					ELSIF TMP_DOUBLE=15 THEN R_COL<="00000100";
					END IF;		
			END CASE;
		ELSIF MOVE=32 THEN
			CASE TMP_DOUBLE IS
					WHEN 0=>R_COL<="00011000";
					WHEN 1=>R_COL<="00011000";
					WHEN 2=>R_COL<="00100100";
					WHEN 3=>R_COL<="00100100";
					WHEN 4=>R_COL<="01000010";
					WHEN 5=>R_COL<="01000010";
					WHEN 6=>R_COL<="10000001";
					WHEN 7=>R_COL<="10000001";
					WHEN 8=>R_COL<="00011000";
					WHEN 9=>R_COL<="00011000";
					WHEN 10=>R_COL<="00100100";
					WHEN 11=>R_COL<="00100100";
					WHEN 12=>R_COL<="01000010";
					WHEN 13=>R_COL<="01000010";
					WHEN 14=>R_COL<="10000001";
					WHEN 15=>R_COL<="10000001";
				END CASE;
		ELSIF MOVE=33 THEN
				IF WIN=1  THEN
					CASE TMP_DOUBLE IS				
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="11000001";
					WHEN 2=>R_COL<="11000001";
					WHEN 3=>R_COL<="11000001";
					WHEN 4=>R_COL<="01111111";
					WHEN 5=>R_COL<="11000001";
					WHEN 6=>R_COL<="11000001";
					WHEN 7=>R_COL<="01111111";
					WHEN 8=>R_COL<="11111111";
					WHEN 9=>R_COL<="11000001";
					WHEN 10=>R_COL<="11000001";
					WHEN 11=>R_COL<="11000001";
					WHEN 12=>R_COL<="01111111";
					WHEN 13=>R_COL<="11000001";
					WHEN 14=>R_COL<="11000001";
					WHEN 15=>R_COL<="01111111";
					END CASE;
				ELSIF WIN=2 THEN
					CASE TMP_DOUBLE IS	
					WHEN 0=>R_COL<="10000001";
					WHEN 1=>R_COL<="01000010";
					WHEN 2=>R_COL<="01000010";
					WHEN 3=>R_COL<="00111100";
					WHEN 4=>R_COL<="00100100";
					WHEN 5=>R_COL<="00011000";
					WHEN 6=>R_COL<="00011000";
					WHEN 7=>R_COL<="00011000";
					WHEN 8=>R_COL<="10000001";
					WHEN 9=>R_COL<="01000010";
					WHEN 10=>R_COL<="01000010";
					WHEN 11=>R_COL<="00111100";
					WHEN 12=>R_COL<="00100100";
					WHEN 13=>R_COL<="00011000";
					WHEN 14=>R_COL<="00011000";
					WHEN 15=>R_COL<="00011000";				
					END CASE;
				ELSE 
					CASE TMP_DOUBLE IS	
					WHEN 0=>R_COL<="10000001";
					WHEN 1=>R_COL<="01000010";
					WHEN 2=>R_COL<="00100100";
					WHEN 3=>R_COL<="00011000";
					WHEN 4=>R_COL<="00011000";
					WHEN 5=>R_COL<="00100100";
					WHEN 6=>R_COL<="01000010";
					WHEN 7=>R_COL<="10000001";
					WHEN 8=>R_COL<="10000001";
					WHEN 9=>R_COL<="01000010";
					WHEN 10=>R_COL<="00100100";
					WHEN 11=>R_COL<="00011000";
					WHEN 12=>R_COL<="00011000";
					WHEN 13=>R_COL<="00100100";
					WHEN 14=>R_COL<="01000010";
					WHEN 15=>R_COL<="10000001";				
					END CASE;
				END IF;
		ELSIF MOVE=0 THEN
			CASE TMP_DOUBLE IS
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="00011000";
					WHEN 2=>R_COL<="00011000";
					WHEN 3=>R_COL<="00011000";
					WHEN 4=>R_COL<="00011000";
					WHEN 5=>R_COL<="00011000";
					WHEN 6=>R_COL<="00011110";
					WHEN 7=>R_COL<="00011000";
					WHEN 8=>R_COL<="11111111";
					WHEN 9=>R_COL<="00011000";
					WHEN 10=>R_COL<="00011000";
					WHEN 11=>R_COL<="00011000";
					WHEN 12=>R_COL<="00011000";
					WHEN 13=>R_COL<="00011000";
					WHEN 14=>R_COL<="00011110";
					WHEN 15=>R_COL<="00011000";
				END CASE;
		ELSIF MOVE=1 THEN
			CASE TMP_DOUBLE IS
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="00000011";
					WHEN 2=>R_COL<="00000011";
					WHEN 3=>R_COL<="00000011";
					WHEN 4=>R_COL<="11111111";
					WHEN 5=>R_COL<="11000000";
					WHEN 6=>R_COL<="11000000";
					WHEN 7=>R_COL<="11111111";
					WHEN 8=>R_COL<="11111111";
					WHEN 9=>R_COL<="00000011";
					WHEN 10=>R_COL<="00000011";
					WHEN 11=>R_COL<="00000011";
					WHEN 12=>R_COL<="11111111";
					WHEN 13=>R_COL<="11000000";
					WHEN 14=>R_COL<="11000000";
					WHEN 15=>R_COL<="11111111";
				END CASE;
		ELSIF MOVE=2 THEN
			CASE TMP_DOUBLE IS
					WHEN 0=>R_COL<="11111111";
					WHEN 1=>R_COL<="10000000";
					WHEN 2=>R_COL<="10000000";
					WHEN 3=>R_COL<="10000000";
					WHEN 4=>R_COL<="11111100";
					WHEN 5=>R_COL<="10000000";
					WHEN 6=>R_COL<="10000000";
					WHEN 7=>R_COL<="11111111";
					WHEN 8=>R_COL<="11111111";
					WHEN 9=>R_COL<="10000000";
					WHEN 10=>R_COL<="10000000";
					WHEN 11=>R_COL<="10000000";
					WHEN 12=>R_COL<="11111100";
					WHEN 13=>R_COL<="10000000";
					WHEN 14=>R_COL<="10000000";
					WHEN 15=>R_COL<="11111111";
				END CASE;	
	END IF;
	END IF;
	END PROCESS;
-------------------------------------------------CHONGZHI
	P12:PROCESS(CLK_ANTISHAKE,RESET_BTN)
		BEGIN
		IF CLK_ANTISHAKE'EVENT AND CLK_ANTISHAKE='1' THEN
		CASE RESET_BTN IS
					WHEN '0'=>RESET<=0;
					WHEN '1'=>RESET<=1;
		END CASE;
	END IF;
	END PROCESS;
-------------------------------------------------SHUMAGUAN
	P13:PROCESS(CLK)
		BEGIN 
		IF CLK'EVENT AND CLK='1' THEN
			IF CAT_TMP=1 THEN 
				CAT_TMP<=0;
			ELSE
				CAT_TMP<=CAT_TMP+1;
			END IF;
		END IF; 
		END PROCESS;
	P14:PROCESS(CLKTMP,MOVE)
	BEGIN
	IF CLKTMP'EVENT AND CLKTMP='1' THEN
		IF MOVE=0 THEN
			MOVE_FLAG<=0;
		ELSIF MOVE=10 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=12 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=14 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=16 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=18 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=20 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=22 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=24 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=26 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=28 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=30 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		ELSIF MOVE=32 THEN
			MOVE_FLAG<=MOVE_FLAG+1;
		END IF;
	END IF;
	END PROCESS;	
	P15:PROCESS(MOVE,CAT_TMP,MOVE_FLAG,CAT_TMP)
		BEGIN
			CASE MOVE IS
			WHEN 0=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
				CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 1=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
				CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 2=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
				CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 3=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 4=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 5=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 6=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 7=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 8=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 9=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 10=>
				NUM_TMP1<="0110000";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 11=>
				NUM_TMP1<="0110000";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 12=>
				NUM_TMP1<="1101101";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 13=>
				NUM_TMP1<="1101101";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 14=>
				NUM_TMP1<="1111001";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 15=>
				NUM_TMP1<="1111001";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 16=>
				NUM_TMP1<="0110011";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 17=>
				NUM_TMP1<="0110011";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 18=>
				NUM_TMP1<="1011011";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 19=>
				NUM_TMP1<="1011011";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 20=>
				NUM_TMP1<="0011111";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 21=>
				NUM_TMP1<="0011111";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 22=>
				NUM_TMP1<="1110000";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 23=>
				NUM_TMP1<="1110000";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 24=>
				NUM_TMP1<="1111111";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 25=>
				NUM_TMP1<="1111111";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 26=>
				NUM_TMP1<="1110011";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 27=>
				NUM_TMP1<="1110011";
				NUM_TMP2<="1111110";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 28=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="0110000";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 29=>
				NUM_TMP1<="1111110";
				NUM_TMP2<="0110000";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 30=>
				NUM_TMP1<="0110000";
				NUM_TMP2<="0110000";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 31=>
				NUM_TMP1<="0110000";
				NUM_TMP2<="0110000";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;
			WHEN 32=>
				NUM_TMP1<="1101101";
				NUM_TMP2<="0110000";
			CASE CAT_TMP IS
				WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
				WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
				END CASE;			
			WHEN 33=>
			CASE MOVE_FLAG IS
				WHEN 0=>
					NUM_TMP1<="1111110";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 1=>
					NUM_TMP1<="0110000";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 2=>
					NUM_TMP1<="1101101";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 3=>
					NUM_TMP1<="1111001";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 4=>
					NUM_TMP1<="0110011";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 5=>
					NUM_TMP1<="1011011";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 6=>
					NUM_TMP1<="0011111";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 7=>
					NUM_TMP1<="1110000";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 8=>
					NUM_TMP1<="1111111";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 9=>
					NUM_TMP1<="1110011";
					NUM_TMP2<="1111110";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 10=>
					NUM_TMP1<="0000001";
					NUM_TMP2<="0110000";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
				WHEN 11=>
					NUM_TMP1<="1101101";
					NUM_TMP2<="0110000";
					CASE CAT_TMP IS				
					WHEN 0=>NUM<=NUM_TMP1;CAT<="11111110";
					WHEN 1=>NUM<=NUM_TMP2;CAT<="11111101";
					END CASE;
			END CASE;
			END CASE;
			
		END PROCESS;
-------------------------------------------------RANDOM
	P16:PROCESS(CLKTMP)
	BEGIN
		IF CLKTMP'EVENT AND CLKTMP='1' THEN
		FEEDBACK<=RAM(3) XNOR RAM(0);
		RAM<=RAM(2 DOWNTO 0)&FEEDBACK;
		END IF;
	END PROCESS;
-------------------------------------------------MULTI
	P17:PROCESS(CLK_ANTISHAKE,MODE_BTN)
		BEGIN
		IF CLK_ANTISHAKE'EVENT AND CLK_ANTISHAKE='1' THEN
		CASE MODE_BTN IS
					WHEN '0'=>MODE_TMP<=0;
					WHEN '1'=>MODE_TMP<=1;
							IF MODE=0 THEN
								MODE<=MODE+1;
							ELSE
								MODE<=0;
							END IF;
		END CASE;
	END IF;
	END PROCESS;
	P18:PROCESS(MODE)
		BEGIN
			IF MODE=0 THEN
				MODE_LIGHT<='1';
			ELSE
				MODE_LIGHT<='0';
			END IF;
		END PROCESS;		
	P19:PROCESS(DTMP)
	BEGIN
		TMP_DOUBLE<=DTMP MOD 16;
	END PROCESS;
	P20:PROCESS(CONTROL_BTN2,CLK_ANTISHAKE)
	BEGIN
	IF CLK_ANTISHAKE'EVENT AND CLK_ANTISHAKE='1' AND FAIL_FLAG=0 THEN
		CASE CONTROL_BTN2 IS
					WHEN "00"=>POSITION2<=POSITION2;
					WHEN "01"=>
						IF POSITION2<7 THEN
							POSITION2<=POSITION2+1;
						END IF;
						
					WHEN "10"=>
						IF POSITION2>0 THEN
							POSITION2<=POSITION2-1;
						END IF;
					WHEN "11"=>POSITION2<=POSITION2;
		END CASE;
	END IF;
	END PROCESS;
-------------------------------------------------LCD
	P21:PROCESS(CLK,NUM_TMP1,NUM_TMP2,MODE,MOVE)
	VARIABLE CNTR:INTEGER RANGE 0 TO 37;
	BEGIN	
			IF CLK'EVENT AND CLK='1' THEN
              CNTR:=CNTR+1;            
          END IF;
          CASE CNTR IS
          -------INIT LCD1602-----------
          WHEN 0 =>RS<='0';QDATA<="00111000";  --0X38,
          WHEN 1 =>RS<='0';QDATA<="00001100";  --0X0C
          WHEN 2 =>RS<='0';QDATA<="00000001";  --0X01
          WHEN 3 =>RS<='0';QDATA<="00000110";  --0X60
          ----------------------------------
          WHEN 4 =>RS<='0';QDATA<="10000000";  --DISPLAY,0X00+0X80,1H1W
          -------DATA DISPLAY-------------
          WHEN 5=>RS<='1';QDATA<="10100000";--�ո�   
		  WHEN 6=>RS<='1';QDATA<="10100000";--�ո�   
		  WHEN 7=>RS<='1';QDATA<="10100000";--�ո�
      WHEN 8=>RS<='1';QDATA<="01001101"; --M   
      WHEN 9=>RS<='1';QDATA<="01001111";--O  
      WHEN 10=>RS<='1';QDATA<="01000100";--D   
      WHEN 11=>RS<='1';QDATA<="01000101";--E   
      WHEN 12=>RS<='1';QDATA<="00111010";--:   
      WHEN 13=>RS<='1';IF MODE=1 THEN QDATA<="01000100";ELSE QDATA<="01010011";END IF;   
      WHEN 14=>RS<='1';IF MODE=1 THEN QDATA<="01001111";ELSE QDATA<="01001001";END IF;     
      WHEN 15=>RS<='1';IF MODE=1 THEN QDATA<="01010101";ELSE QDATA<="01001110";END IF;   
      WHEN 16=>RS<='1';IF MODE=1 THEN QDATA<="01000010";ELSE QDATA<="01000111";END IF;   
      WHEN 17=>RS<='1';IF MODE=1 THEN QDATA<="01001100";ELSE QDATA<="01001100";END IF;  
      WHEN 18=>RS<='1';IF MODE=1 THEN QDATA<="01000101";ELSE QDATA<="01000101";END IF;   
      WHEN 19=>RS<='1';QDATA<="10100000";---�ո�   
      WHEN 20=>RS<='1';QDATA<="10100000";---�ո�
     ---------------------------
        WHEN 21=>RS<='0';QDATA<="11000000";--�趨��ʾ��λ����10H+80H��
       ----------------------------
       WHEN 22=>RS<='1';QDATA<="10100000";---�ո�   
     WHEN 23=>RS<='1';QDATA<="10100000";---�ո�   
     WHEN 24=>RS<='1';QDATA<="10100000";---�ո�  
     WHEN 25=>RS<='1';QDATA<="01010011";---S  
     WHEN 26=>RS<='1';QDATA<="01000011";---C   
     WHEN 27=>RS<='1';QDATA<="01001111";---O
     WHEN 28=>RS<='1';QDATA<="01010010";--R   
     WHEN 29=>RS<='1';QDATA<="01000101";---E   
     WHEN 30=>RS<='1';QDATA<="00111010";---:   
     WHEN 31=>RS<='1';
			IF NUM_TMP2="0110000" THEN QDATA<="00110001";
			ELSIF NUM_TMP2="1111110" THEN QDATA<="00110000";
			END IF;
     WHEN 32=>RS<='1';
			IF NUM_TMP1="1111110" THEN QDATA<="00110000";
			ELSIF NUM_TMP1="0110000" THEN QDATA<="00110001";
			ELSIF NUM_TMP1="1101101" THEN QDATA<="00110010";
			ELSIF NUM_TMP1="1111001" THEN QDATA<="00110011";
			ELSIF NUM_TMP1="0110011" THEN QDATA<="00110100";
			ELSIF NUM_TMP1="1011011" THEN QDATA<="00110101";
			ELSIF NUM_TMP1="0011111" THEN QDATA<="00110110";
			ELSIF NUM_TMP1="1110000" THEN QDATA<="00110111";
			ELSIF NUM_TMP1="1111111" THEN QDATA<="00111000";
			ELSIF NUM_TMP1="1110011" THEN QDATA<="00111001";
			
			END IF;
     WHEN 33=>RS<='1';QDATA<="10100000";---�ո�  
     WHEN 34=>RS<='1';QDATA<="10100000";---�ո� 
     WHEN 35=>RS<='1';QDATA<="10100000";---�ո� 
     WHEN 36=>RS<='1';QDATA<="10100000";---�ո� 
     WHEN 37=>RS<='1';QDATA<="10100000";---�ո� 
     END CASE;
	END PROCESS;
-------------------------------------------------MUSIC
	P22:PROCESS(CLK_IN)
		BEGIN
			IF CLK_IN'EVENT AND CLK_IN='1' THEN
				IF TMP_SOUND=6249999 THEN
					TMP_SOUND<=0;
					CLK_SOUND<=NOT CLK_SOUND;
				ELSE
					TMP_SOUND<=TMP_SOUND+1;
				END IF;
			END IF;			
		END PROCESS;
	P23:PROCESS(CLK_SOUND)
		BEGIN
			IF CLK_SOUND'EVENT AND CLK_SOUND='1'THEN
				IF SELECTION=127 THEN
					SELECTION<=0;
				ELSE
					SELECTION<=SELECTION+1;
				END IF;
			END IF;
			CASE SELECTION IS
			WHEN 0=>TUNE<=MI;
			WHEN 1=>TUNE<=FA;
			WHEN 2=>TUNE<=SO;
			WHEN 3=>TUNE<=SO;
			WHEN 4=>TUNE<=MI;
			WHEN 5=>TUNE<=MI;
			WHEN 6=>TUNE<=XI;
			WHEN 7=>TUNE<=0;
			WHEN 8=>TUNE<=MI;
			WHEN 9=>TUNE<=FA;
			WHEN 10=>TUNE<=SO;
			WHEN 11=>TUNE<=SO;
			WHEN 12=>TUNE<=MI;
			WHEN 13=>TUNE<=MI;
			WHEN 14=>TUNE<=XI;
			WHEN 15=>TUNE<=XI;
			WHEN 16=>TUNE<=0;
			WHEN 17=>TUNE<=0;
			WHEN 18=>TUNE<=XI;
			WHEN 19=>TUNE<=DO_HIGH;
			WHEN 20=>TUNE<=XI;
			WHEN 21=>TUNE<=LA;
			WHEN 22=>TUNE<=SO;
			WHEN 23=>TUNE<=0;
			WHEN 24=>TUNE<=SO;
			WHEN 25=>TUNE<=FA;
			WHEN 26=>TUNE<=MI;
			WHEN 27=>TUNE<=MI;
			WHEN 28=>TUNE<=0;
			WHEN 29=>TUNE<=0;
			WHEN 30=>TUNE<=0;
			WHEN 31=>TUNE<=0;
			WHEN 32=>TUNE<=MI;
			WHEN 33=>TUNE<=FA;
			WHEN 34=>TUNE<=SO;
			WHEN 35=>TUNE<=SO;
			WHEN 36=>TUNE<=MI;
			WHEN 37=>TUNE<=MI;
			WHEN 38=>TUNE<=0;
			WHEN 39=>TUNE<=0;
			
			WHEN 40=>TUNE<=SO;
			WHEN 41=>TUNE<=LA;
			WHEN 42=>TUNE<=XI;
			WHEN 43=>TUNE<=XI;
			WHEN 44=>TUNE<=MI;
			WHEN 45=>TUNE<=MI;
			WHEN 46=>TUNE<=0;
			WHEN 47=>TUNE<=0;
			
			WHEN 48=>TUNE<=RE_HIGH;
			WHEN 49=>TUNE<=DO_HIGH2;
			WHEN 50=>TUNE<=RE_HIGH;
			WHEN 51=>TUNE<=DO_HIGH2;
			WHEN 52=>TUNE<=RE_HIGH;
			WHEN 53=>TUNE<=DO_HIGH2;
			WHEN 54=>TUNE<=RE_HIGH;
			WHEN 55=>TUNE<=MI_HIGH;
			WHEN 56=>TUNE<=RE_HIGH;
			WHEN 57=>TUNE<=DO_HIGH2;
			WHEN 58=>TUNE<=XI;
			WHEN 59=>TUNE<=XI;
			WHEN 60=>TUNE<=0;
			WHEN 61=>TUNE<=0;
			WHEN 62=>TUNE<=0;
			WHEN 63=>TUNE<=0;
			WHEN 64=>TUNE<=XI;
			WHEN 65=>TUNE<=DO_HIGH2;
			WHEN 66=>TUNE<=RE_HIGH;
			WHEN 67=>TUNE<=0;
			WHEN 68=>TUNE<=RE_HIGH;
			WHEN 69=>TUNE<=0;
			WHEN 70=>TUNE<=RE_HIGH;
			WHEN 71=>TUNE<=0;
			WHEN 72=>TUNE<=RE_HIGH;
			WHEN 73=>TUNE<=0;
			WHEN 74=>TUNE<=RE_HIGH;
			WHEN 75=>TUNE<=MI_HIGH;
			WHEN 76=>TUNE<=RE_HIGH;
			WHEN 77=>TUNE<=DO_HIGH2;
			WHEN 78=>TUNE<=RE_HIGH;
			WHEN 79=>TUNE<=0;
			WHEN 80=>TUNE<=XI;
			WHEN 81=>TUNE<=DO_HIGH2;
			WHEN 82=>TUNE<=RE_HIGH;
			WHEN 83=>TUNE<=0;
			WHEN 84=>TUNE<=RE_HIGH;
			WHEN 85=>TUNE<=0;	
			WHEN 86=>TUNE<=RE_HIGH;
			WHEN 87=>TUNE<=0;	
			WHEN 88=>TUNE<=RE_HIGH;
			WHEN 89=>TUNE<=DO_HIGH2;
			WHEN 90=>TUNE<=XI;
			WHEN 91=>TUNE<=XI;
			WHEN 92=>TUNE<=0;
			WHEN 93=>TUNE<=0;	
			WHEN 94=>TUNE<=0;
			WHEN 95=>TUNE<=0;
			WHEN 96=>TUNE<=XI;
			WHEN 97=>TUNE<=DO_HIGH2;
			WHEN 98=>TUNE<=RE_HIGH;
			WHEN 99=>TUNE<=0;
			WHEN 100=>TUNE<=RE_HIGH;
			WHEN 101=>TUNE<=0;
			WHEN 102=>TUNE<=RE_HIGH;
			WHEN 103=>TUNE<=0;
			WHEN 104=>TUNE<=RE_HIGH;
			WHEN 105=>TUNE<=0;
			WHEN 106=>TUNE<=RE_HIGH;
			WHEN 107=>TUNE<=MI_HIGH;
			WHEN 108=>TUNE<=RE_HIGH;
			WHEN 109=>TUNE<=DO_HIGH2;
			WHEN 110=>TUNE<=RE_HIGH;
			WHEN 111=>TUNE<=0;
			WHEN 112=>TUNE<=XI;
			WHEN 113=>TUNE<=DO_HIGH2;
			WHEN 114=>TUNE<=RE_HIGH;
			WHEN 115=>TUNE<=0;
			WHEN 116=>TUNE<=RE_HIGH;
			WHEN 117=>TUNE<=0;	
			WHEN 118=>TUNE<=RE_HIGH;
			WHEN 119=>TUNE<=0;	
			WHEN 120=>TUNE<=RE_HIGH;
			WHEN 121=>TUNE<=DO_HIGH2;
			WHEN 122=>TUNE<=XI;
			WHEN 123=>TUNE<=XI;	
			WHEN 124=>TUNE<=0;
			WHEN 125=>TUNE<=0;	
			WHEN 126=>TUNE<=0;
			WHEN 127=>TUNE<=0;		
			END CASE;
			
		END PROCESS;	
	P24:PROCESS(CLK_IN,TUNE)
		BEGIN
			IF CLK_IN'EVENT AND CLK_IN='1'THEN
				IF CNT=TUNE OR CNT>TUNE THEN
					CNT<=0;
					CLK_BEEP<=NOT CLK_BEEP;
				ELSE
					CNT<=CNT+1;
				END IF;
			END IF;
			BEEP<=CLK_BEEP;
		END PROCESS;	
END IGNIGHT;